package types;
    typedef logic [31:0] word_t;
endpackage
