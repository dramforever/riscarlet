package rscl_types;
    typedef logic [31:0]    word_t;
    typedef logic [3:0]     bsel_t;

    typedef logic [31:0]    instr_t;
    typedef logic [4:0]     rnum_t;
    typedef logic [6:0]     opcode_t;
    typedef logic [6:0]     funct7_t;
    typedef logic [2:0]     funct3_t;

    typedef logic [3:0]     cause_t;
    typedef logic [11:0]    csr_num_t;
endpackage
