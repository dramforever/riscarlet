`include "prim/multiply_signed.sv"
`include "prim/multiply.sv"
