`include "riscv/types.sv"

`include "wishbone/wishbone.sv"
`include "riscv/pipeline.sv"
`include "riscv/regport.sv"

`include "riscv/riscv_alu.sv"

`include "riscv/pipe_slice.sv"
`include "riscv/stage_fetch.sv"
`include "riscv/riscarlet.sv"
