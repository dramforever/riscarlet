`include "riscv/types.sv"

`include "bus/bus.sv"
`include "bus/bus_req_c.sv"
`include "bus/bus_rsp_c.sv"
`include "riscv/pipeline.sv"
`include "riscv/regport.sv"

`include "riscv/riscv_alu.sv"

`include "riscv/pipe_slice.sv"
`include "riscv/stage_fetch.sv"
`include "riscv/riscarlet.sv"
