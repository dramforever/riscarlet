module rscl_top();
endmodule
